*Tamrin1ForMinTerm
.INCLUDE	model.txt

*===>NAME	+	-	VALUE
VCC VCC 0 5
*===>NAME	+	-	PULSE(MIN MAX DELAYTIME RISETIME FALLTIME PULSEWIDTH DORETANAVON)
VIN	IN 	0		PULSE(0 5 0N 10N 10N 200N 500N)
R1	IN	OUTR1	10K
*==>TRANZISTOR BYPOLAR => QNAME	  COLLECTOR  	BASE   EMMITER  NPN
Q1	OUT OUTR1 	0 NPN
R2	VCC OUT   	1K
*=>.DC	iNPUT	START	STOP	STEP 	MEHVAR_OFOGHI	
.DC	VG	0		5	0.1
*=> .PRINT DC V(1) I(5)=>MEHVAR AMOODI NESBAT BE DC
*=> mEVAR OFOGHI TIME BASHE .TRAN	200P	20N		(START = 10NS)


